module 4_to_16_encoder (
    ports
);
    
endmodule