library verilog;
use verilog.vl_types.all;
entity phase3_tb is
end phase3_tb;
