module  sub_32_bit (
    input [31:0] 
);
//to subtract, you need to negate the second number, then add it to first
//To negate a number, you need the two's compliment, which is done by
//taking the inverse of the number, then adding 1 to it.
    
endmodule