module multiplication_32_bit (
  input [31:0] a, b,
  output [31:0] hi, lo,

);
  
endmodule