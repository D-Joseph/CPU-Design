module selectencodelogic (
    input [31:0] instruction,
    input Gra, Grb, Grc, Rin, Rout, BAout,
    output [31:0] C_Sign_Extended,
    output [15:0] RegIn, RegOut,
    
);
    
endmodule